module c ();
  d u_d();
endmodule
