module a ();
  b u_b();
  c u_c();
endmodule
