module b ();
  c u_c();
endmodule
