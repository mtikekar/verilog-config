module d ();
endmodule
